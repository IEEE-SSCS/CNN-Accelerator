module img2col(
    
);
    





endmodule