module parameter_calc(
    input logic stride , input logic 
);
    

always_comb begin
    



end

endmodule